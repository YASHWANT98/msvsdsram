// Generated for: spectre
// Generated on: May 10 08:51:04 2023
// Design library name: SCL180_Design
// Design cell name: 1_bit_SRAM
// Design view name: schematic
simulator lang=spectre
global 0

// Library name: SCL180_Design
// Cell name: 1_bit_SRAM
// View name: schematic
M27 (Out BL net65 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M26 (net66 BLbar net65 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M25 (Dout Out 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M24 (net65 Rd_EN 0 0) n18 w=1.26 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M19 (net70 Vin 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M18 (net67 net70 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M12 (net68 net67 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M11 (net68 WR_EN 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M16 (net71 net70 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M15 (net71 WR_EN 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M14 (0 net71 BLbar 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M13 (0 net68 BL 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M2 (BL WL BL 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 m=1
M3 (BLbar WL BLbar 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M0 (BLbar BL 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M1 (BL BLbar 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M30 (net66 net66 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M29 (Dout Out VDD VDD) p18 w=0.84 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M28 (Out net66 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M23 (BL Precharge VDD VDD) p18 w=0.84 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M22 (BLbar Precharge VDD VDD) p18 w=0.84 l=0.18 as=0.1984 ad=0.1984 \
        ps=1.88 pd=1.88 m=1
M21 (net67 net70 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M20 (net70 Vin VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M17 (net69 net67 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M10 (net68 WR_EN net69 VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M9 (VDD net70 net72 VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M8 (net72 WR_EN net71 VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M7 (BLbar 0 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M6 (VDD 0 BL VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M5 (BL BLbar VDD VDD) p18 w=0.84 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M4 (BLbar BL VDD VDD) p18 w=0.84 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
V2 (Rd_EN 0) vsource type=pulse val0=1.8 val1=0 period=10n width=5n
V1 (Precharge 0) vsource type=pulse val0=0 val1=1.8 period=10n width=5n
V0 (VDD 0) vsource dc=1.8 type=dc
simulatorOptions options psfversion="1.4.0" reltol=1e-3 vabstol=1e-6 \
    iabstol=1e-12 temp=27 tnom=27 scalem=1.0 scale=1.0 gmin=1e-12 rforce=1 \
    maxnotes=5 maxwarns=5 digits=5 cols=80 pivrel=1e-3 \
    sensfile="../psf/sens.output" checklimitdest=psf 
modelParameter info what=models where=rawfile
element info what=inst where=rawfile
outputParameter info what=output where=rawfile
designParamVals info what=parameters where=rawfile
primitives info what=primitives where=rawfile
subckts info what=subckts where=rawfile
saveOptions options save=allpub
