// Generated for: spectre
// Generated on: May 10 06:34:39 2023
// Design library name: SCL180_Design
// Design cell name: D_flipflop
// Design view name: schematic
simulator lang=spectre
global 0

// Library name: SCL180_Design
// Cell name: D_flipflop
// View name: schematic
M17 (net1 CLK net4 net4) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M7 (VDD Q net4 VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M6 (Q net1 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M5 (net3 CLKbar net1 net3) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M4 (net3 net6 VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M3 (CLKbar CLK VDD VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M2 (VDD net3 net2 VDD) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M1 (net6 CLKbar net2 net2) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M0 (D CLK net6 D) p18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M16 (net1 CLKbar net4 net4) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M15 (0 Q net4 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 m=1
M14 (Q net1 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 m=1
M13 (net3 CLK net1 net3) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M12 (net3 net6 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M11 (CLKbar CLK 0 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M10 (0 net3 net2 0) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
M9 (net6 CLK net2 net2) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 \
        pd=1.88 m=1
M8 (D CLKbar net6 D) n18 w=0.42 l=0.18 as=0.1984 ad=0.1984 ps=1.88 pd=1.88 \
        m=1
V0 (VDD 0) vsource dc=1.8 type=dc
V2 (D 0) vsource type=pulse val0=0 val1=1.8 period=30n delay=2.5n \
        width=15n
V1 (CLK 0) vsource type=pulse val0=1.8 val1=0 period=10n width=5n
simulatorOptions options psfversion="1.4.0" reltol=1e-3 vabstol=1e-6 \
    iabstol=1e-12 temp=27 tnom=27 scalem=1.0 scale=1.0 gmin=1e-12 rforce=1 \
    maxnotes=5 maxwarns=5 digits=5 cols=80 pivrel=1e-3 \
    sensfile="../psf/sens.output" checklimitdest=psf 
modelParameter info what=models where=rawfile
element info what=inst where=rawfile
outputParameter info what=output where=rawfile
designParamVals info what=parameters where=rawfile
primitives info what=primitives where=rawfile
subckts info what=subckts where=rawfile
saveOptions options save=allpub
